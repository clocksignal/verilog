//module Half_Adder(
//        input [1:0] IN,
//        output [1:0] OUT
//    );
    
//    wire A = IN[0];
//    wire B = IN[1];
//    // SUM
//    xor(OUT[0],A,B);
//    // Carry out
//    and(OUT[1],A,B);
//endmodule
