module barrel_shifter_12bits(
        input [11:0]IN,
        input [1:0] select,
        output [11:0] OUT
    );
    //barrel_shifter UUT1(.IN({IN[3],IN[2],IN[1],IN[0]}),.select(),.OUT());
    
endmodule
